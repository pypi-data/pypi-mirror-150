//
//  ITC99 Benchmark
//  Downloaded from http://www.cad.polito.it/tools/itc99.html
//  
//  ----------------------------------------------------------------------
//  
//  This netlist was generated with Cadence RTL Compiler in a quick 
//  synthesis run.
//  
//  ----------------------------------------------------------------------
//  
//  Copyright (C) 1999
//  Fulvio Corno, Matteo Sonze Reorda, Giovanni Squillero
//  Politecnico di Torino
//  
//  This source file may be used and distributed without restriction
//  provided that this copyright statement is not removed from the
//  file and that any derivative work contains the original copyright
//  notice and the associated disclaimer.
//  
//  This source file is free software; you can redistribute it and/or
//  modify it under the terms of the GNU General Public License as
//  published by the Free Software Foundation.
//  
//  This source is distributed in the hope that it will be useful,
//  but WITHOUT ANY WARRANTY; without even the implied warranty of
//  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
//  General Public License for more details.
//  
//  You should have received a copy of the GNU General Public License
//  along with this source; if not, download it from
//  http://www.gnu.org/copyleft/gpl.html
//  

// Generated by Cadence RTL Compiler (RC) v05.10-b006_1

module b10(r_button, g_button, key, start, reset, test, cts, ctr, rts,
     rtr, clock, v_in, v_out);
  input r_button, g_button, key, start, reset, test, rts, rtr, clock;
  input [3:0] v_in;
  output cts, ctr;
  output [3:0] v_out;
  wire r_button, g_button, key, start, reset, test, rts, rtr, clock;
  wire [3:0] v_in;
  wire cts, ctr;
  wire [3:0] v_out;
  wire n_1, n_2, n_4, n_5, n_6, n_7, n_8, n_9;
  wire n_12, n_13, n_15, n_16, n_17, n_18, n_20, n_21;
  wire n_22, n_24, n_27, n_29, n_30, n_31, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_45, n_46, n_47;
  wire n_49, n_57, n_59, n_60, n_61, n_63, n_67, n_72;
  wire n_73, n_74, n_75, n_77, n_78, n_79, n_80, n_85;
  wire n_86, n_87, n_89, n_90, n_91, n_92, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_103, n_104, n_110, n_111;
  wire n_112, n_113, n_115, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_131, n_132, n_133, n_135;
  wire n_137, n_138, n_140, n_141, n_142, n_145, n_148, n_149;
  wire n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_161;
  wire n_162, n_163, n_165, n_166, n_167, n_168, n_169, n_171;
  wire n_174, n_175, n_176, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_186, n_188, n_189, n_190, n_191, n_192;
  wire n_194, n_195, n_196, n_197, n_199, n_200, n_201, n_203;
  wire n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211;
  wire n_212, n_213, n_214, n_215, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_233, n_235, n_238, n_241, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261;
  wire n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269;
  wire n_270, n_271, n_274, n_276, n_277, n_279, n_280, n_281;
  wire n_282, n_284, n_285, n_286, n_287, n_288, n_289, n_292;
  wire n_293, n_294, n_295, n_297, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_307, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_322;
  wire n_323, n_324, n_325, n_328, n_329, n_330, n_331, n_332;
  wire n_333, n_335, n_336, n_337, n_338, n_339, n_340, n_348;
  wire n_350, n_351, n_352, n_358, n_377, n_381, n_388, n_389;
  wire n_391, n_392, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_411;
  wire n_412, n_413, n_414, n_415, n_416, n_430, n_431, n_432;
  wire n_433, n_441, n_442, n_443, n_444, n_445, n_446, n_447;
  wire n_449, n_451, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, stato, stato_5, stato_6, stato_7;
  wire voto2;
  DFFSRX1 \stato_reg[2] (.RN (n_340), .SN (1'b1), .CK (clock), .D
       (n_339), .Q (stato_6), .QN ());
  DFFSRX1 \stato_reg[0] (.RN (n_340), .SN (1'b1), .CK (clock), .D
       (n_446), .Q (stato), .QN ());
  DFFSRX1 voto1_reg(.RN (n_340), .SN (1'b1), .CK (clock), .D (n_336),
       .Q (n_178), .QN ());
  DFFSRX1 \stato_reg[1] (.RN (n_340), .SN (1'b1), .CK (clock), .D
       (n_333), .Q (stato_5), .QN ());
  DFFSRX1 \v_out_reg[2] (.RN (n_340), .SN (1'b1), .CK (clock), .D
       (n_337), .Q (v_out[2]), .QN ());
  DFFSRX1 \v_out_reg[3] (.RN (n_340), .SN (1'b1), .CK (clock), .D
       (n_332), .Q (v_out[3]), .QN ());
  DFFSRX1 cts_reg(.RN (n_340), .SN (1'b1), .CK (clock), .D (n_335), .Q
       (cts), .QN ());
  DFFSRX1 \v_out_reg[0] (.RN (n_340), .SN (1'b1), .CK (clock), .D
       (n_331), .Q (v_out[0]), .QN ());
  DFFSRX1 \v_out_reg[1] (.RN (n_340), .SN (1'b1), .CK (clock), .D
       (n_338), .Q (v_out[1]), .QN ());
  OR4X1 g1181(.A (n_189), .B (n_238), .C (n_195), .D (n_324), .Y
       (n_339));
  DFFSRX1 last_g_reg(.RN (n_340), .SN (1'b1), .CK (clock), .D (n_330),
       .Q (n_300), .QN ());
  DFFSRX1 last_r_reg(.RN (n_340), .SN (1'b1), .CK (clock), .D (n_329),
       .Q (n_38), .QN ());
  DFFSRX1 \sign_reg[3] (.RN (n_340), .SN (1'b1), .CK (clock), .D
       (n_328), .Q (n_286), .QN ());
  DFFSRX1 ctr_reg(.RN (n_340), .SN (1'b1), .CK (clock), .D (n_416), .Q
       (ctr), .QN ());
  NAND2X2 g1210(.A (n_316), .B (n_260), .Y (n_338));
  NAND2X2 g1211(.A (n_315), .B (n_264), .Y (n_337));
  DFFSRX1 voto2_reg(.RN (n_340), .SN (1'b1), .CK (clock), .D (n_325),
       .Q (voto2), .QN ());
  DFFSRX1 \stato_reg[3] (.RN (n_340), .SN (1'b1), .CK (clock), .D
       (n_323), .Q (stato_7), .QN ());
  NAND2X1 g1199(.A (n_467), .B (n_468), .Y (n_336));
  NAND3X1 g1216(.A (n_313), .B (n_254), .C (n_271), .Y (n_335));
  NAND3X1 g1202(.A (n_322), .B (n_305), .C (n_209), .Y (n_333));
  NAND2X2 g1205(.A (n_320), .B (n_263), .Y (n_332));
  NAND2X2 g1209(.A (n_319), .B (n_261), .Y (n_331));
  DFFSRX1 voto3_reg(.RN (n_340), .SN (1'b1), .CK (clock), .D (n_309),
       .Q (n_27), .QN ());
  NAND3X1 g1217(.A (n_312), .B (n_301), .C (n_225), .Y (n_330));
  NAND3X1 g1218(.A (n_311), .B (n_279), .C (n_222), .Y (n_329));
  NAND2X1 g1208(.A (n_351), .B (n_352), .Y (n_328));
  DFFSRX1 voto0_reg(.RN (n_340), .SN (1'b1), .CK (clock), .D (n_302),
       .Q (n_47), .QN ());
  NAND4X1 g1200(.A (n_274), .B (n_250), .C (n_281), .D (n_282), .Y
       (n_325));
  OAI21X1 g1214(.A0 (n_196), .A1 (n_74), .B0 (n_297), .Y (n_324));
  NAND4X1 g1201(.A (n_247), .B (n_205), .C (n_303), .D (n_265), .Y
       (n_323));
  AOI21X1 g1221(.A0 (n_86), .A1 (n_175), .B0 (n_304), .Y (n_322));
  INVX1 g1203(.A (n_307), .Y (n_467));
  AOI22X1 g1231(.A0 (n_318), .A1 (v_out[3]), .B0 (n_317), .B1
       (v_out[3]), .Y (n_320));
  AOI22X1 g1232(.A0 (n_318), .A1 (v_out[0]), .B0 (n_317), .B1
       (v_out[0]), .Y (n_319));
  AOI22X1 g1233(.A0 (n_314), .A1 (v_out[1]), .B0 (n_317), .B1
       (v_out[1]), .Y (n_316));
  AOI22X1 g1234(.A0 (n_314), .A1 (v_out[2]), .B0 (n_317), .B1
       (v_out[2]), .Y (n_315));
  AOI22X1 g1235(.A0 (n_433), .A1 (cts), .B0 (n_169), .B1 (cts), .Y
       (n_313));
  OAI21X1 g1237(.A0 (n_258), .A1 (n_310), .B0 (n_300), .Y (n_312));
  OAI21X1 g1238(.A0 (n_257), .A1 (n_310), .B0 (n_38), .Y (n_311));
  NAND3X1 g1212(.A (n_289), .B (n_268), .C (n_267), .Y (n_309));
  AOI22X1 g1247(.A0 (n_255), .A1 (n_286), .B0 (n_358), .B1 (n_286), .Y
       (n_352));
  NAND4X1 g1204(.A (n_252), .B (n_284), .C (n_231), .D (n_245), .Y
       (n_307));
  NOR2X1 g1227(.A (n_288), .B (n_285), .Y (n_351));
  AOI21X1 g1230(.A0 (n_407), .A1 (n_269), .B0 (n_295), .Y (n_305));
  NAND2X1 g1245(.A (n_270), .B (n_303), .Y (n_304));
  NAND4X1 g1219(.A (n_277), .B (n_201), .C (n_233), .D (n_211), .Y
       (n_302));
  NAND2X1 g1264(.A (n_259), .B (n_300), .Y (n_301));
  NOR2X1 g1226(.A (n_243), .B (n_280), .Y (n_297));
  NAND3X1 g1236(.A (n_469), .B (n_194), .C (n_294), .Y (n_295));
  NAND2X1 g1257(.A (n_293), .B (n_292), .Y (n_318));
  NAND2X1 g1259(.A (n_293), .B (n_292), .Y (n_314));
  AOI22X1 g1229(.A0 (n_276), .A1 (n_27), .B0 (n_112), .B1 (n_251), .Y
       (n_289));
  AND2X1 g1294(.A (n_287), .B (n_286), .Y (n_288));
  OAI21X1 g1240(.A0 (n_181), .A1 (n_18), .B0 (n_149), .Y (n_285));
  INVX1 g1241(.A (n_248), .Y (n_284));
  AOI21X1 g1243(.A0 (n_59), .A1 (n_407), .B0 (n_213), .Y (n_282));
  AOI21X1 g1244(.A0 (n_266), .A1 (voto2), .B0 (n_208), .Y (n_281));
  NAND4X1 g1246(.A (n_165), .B (n_294), .C (n_162), .D (n_152), .Y
       (n_280));
  OAI21X1 g1250(.A0 (n_226), .A1 (n_453), .B0 (n_38), .Y (n_279));
  NAND2X1 g1251(.A (n_276), .B (n_47), .Y (n_277));
  NAND2X1 g1253(.A (n_276), .B (n_244), .Y (n_468));
  NAND2X1 g1255(.A (n_276), .B (voto2), .Y (n_274));
  OAI21X1 g1262(.A0 (n_317), .A1 (n_407), .B0 (cts), .Y (n_271));
  NAND2X1 g1265(.A (n_203), .B (n_269), .Y (n_270));
  AOI21X1 g1266(.A0 (n_89), .A1 (n_249), .B0 (n_408), .Y (n_268));
  AOI21X1 g1268(.A0 (n_266), .A1 (n_27), .B0 (n_229), .Y (n_267));
  AOI21X1 g1269(.A0 (n_230), .A1 (n_154), .B0 (n_235), .Y (n_265));
  AOI21X1 g1271(.A0 (n_262), .A1 (v_out[2]), .B0 (n_228), .Y (n_264));
  AOI21X1 g1272(.A0 (n_262), .A1 (v_out[3]), .B0 (n_224), .Y (n_263));
  AOI21X1 g1273(.A0 (n_262), .A1 (v_out[0]), .B0 (n_220), .Y (n_261));
  AOI21X1 g1274(.A0 (n_262), .A1 (v_out[1]), .B0 (n_219), .Y (n_260));
  NAND2X1 g1277(.A (n_292), .B (n_392), .Y (n_259));
  NAND2X1 g1285(.A (n_227), .B (n_256), .Y (n_258));
  NAND2X1 g1290(.A (n_292), .B (n_256), .Y (n_257));
  NAND2X1 g1293(.A (n_207), .B (n_292), .Y (n_255));
  AOI21X1 g1300(.A0 (rtr), .A1 (n_175), .B0 (n_192), .Y (n_254));
  AOI22X1 g1303(.A0 (n_249), .A1 (n_90), .B0 (n_251), .B1 (n_178), .Y
       (n_252));
  AOI22X1 g1304(.A0 (n_249), .A1 (n_80), .B0 (n_251), .B1 (voto2), .Y
       (n_250));
  OAI21X1 g1242(.A0 (n_212), .A1 (n_127), .B0 (n_167), .Y (n_248));
  AOI21X1 g1215(.A0 (n_171), .A1 (n_246), .B0 (n_184), .Y (n_247));
  NAND2X1 g1329(.A (n_389), .B (n_191), .Y (n_287));
  NAND2X1 g1254(.A (n_183), .B (n_244), .Y (n_245));
  NAND2X1 g1352(.A (n_389), .B (n_432), .Y (n_243));
  INVX1 g1224(.A (n_210), .Y (n_241));
  INVX1 g1288(.A (n_206), .Y (n_238));
  NOR2X1 g1292(.A (n_453), .B (n_358), .Y (n_293));
  OAI21X1 g1298(.A0 (n_256), .A1 (test), .B0 (n_168), .Y (n_235));
  NAND2X1 g1299(.A (n_166), .B (n_269), .Y (n_469));
  AOI22X1 g1301(.A0 (n_249), .A1 (n_94), .B0 (n_47), .B1 (n_460), .Y
       (n_233));
  AOI21X1 g1302(.A0 (n_230), .A1 (v_in[1]), .B0 (n_179), .Y (n_231));
  OAI21X1 g1306(.A0 (n_215), .A1 (n_6), .B0 (n_176), .Y (n_229));
  NOR2X1 g1312(.A (n_78), .B (n_223), .Y (n_228));
  OR2X1 g1319(.A (n_186), .B (n_175), .Y (n_310));
  INVX1 g1322(.A (n_226), .Y (n_227));
  INVX4 g1324(.A (n_199), .Y (n_292));
  AOI22X1 g1248(.A0 (n_121), .A1 (n_407), .B0 (n_300), .B1 (n_221), .Y
       (n_225));
  NOR2X1 g1332(.A (n_95), .B (n_223), .Y (n_224));
  AOI22X1 g1249(.A0 (n_120), .A1 (n_407), .B0 (n_38), .B1 (n_221), .Y
       (n_222));
  NOR2X1 g1341(.A (n_96), .B (n_223), .Y (n_220));
  NOR2X1 g1344(.A (n_92), .B (n_223), .Y (n_219));
  NAND2X1 g1256(.A (n_156), .B (n_72), .Y (n_218));
  AOI21X1 g1220(.A0 (n_111), .A1 (n_188), .B0 (n_223), .Y (n_214));
  NOR2X1 g1263(.A (n_124), .B (n_212), .Y (n_213));
  AOI22X1 g1270(.A0 (n_153), .A1 (n_47), .B0 (n_18), .B1 (n_221), .Y
       (n_211));
  NAND4X1 g1225(.A (n_209), .B (n_138), .C (n_131), .D (n_126), .Y
       (n_210));
  OAI21X1 g1275(.A0 (n_182), .A1 (n_79), .B0 (n_180), .Y (n_208));
  NAND2X2 g1279(.A (n_207), .B (n_191), .Y (n_276));
  NAND3X1 g1289(.A (rtr), .B (n_204), .C (n_163), .Y (n_206));
  NAND3X1 g1291(.A (rtr), .B (n_204), .C (n_154), .Y (n_205));
  NAND2X1 g1296(.A (n_215), .B (n_377), .Y (n_203));
  AOI22X1 g1305(.A0 (n_230), .A1 (v_in[0]), .B0 (n_91), .B1 (n_409), .Y
       (n_201));
  NAND2X1 g1310(.A (n_407), .B (n_72), .Y (n_200));
  NAND2X1 g1318(.A (n_256), .B (n_432), .Y (n_262));
  NAND2X1 g1323(.A (n_123), .B (n_190), .Y (n_226));
  NAND2X2 g1325(.A (n_148), .B (n_145), .Y (n_199));
  NAND2X1 g1334(.A (n_432), .B (n_457), .Y (n_266));
  NAND2X1 g1335(.A (n_161), .B (n_196), .Y (n_197));
  INVX1 g1338(.A (n_194), .Y (n_195));
  NAND2X1 g1342(.A (n_141), .B (n_133), .Y (n_358));
  NOR2X1 g1347(.A (n_20), .B (n_191), .Y (n_192));
  NAND2X1 g1349(.A (n_388), .B (n_190), .Y (n_317));
  AOI21X1 g1222(.A0 (n_75), .A1 (n_188), .B0 (n_191), .Y (n_189));
  NOR2X1 g1223(.A (n_155), .B (n_191), .Y (n_184));
  NAND2X1 g1281(.A (n_182), .B (n_432), .Y (n_183));
  AOI21X1 g1295(.A0 (test), .A1 (n_132), .B0 (n_221), .Y (n_181));
  NAND2X1 g1309(.A (n_230), .B (v_in[2]), .Y (n_180));
  NAND3X1 g1311(.A (start), .B (n_122), .C (n_140), .Y (n_212));
  AND2X1 g1313(.A (n_178), .B (n_460), .Y (n_179));
  NAND2X1 g1314(.A (n_175), .B (n_398), .Y (n_176));
  NOR2X1 g1315(.A (n_196), .B (n_99), .Y (n_174));
  NAND2X1 g1320(.A (n_406), .B (n_1), .Y (n_209));
  NAND2X1 g1326(.A (n_230), .B (n_103), .Y (n_303));
  NOR2X1 g1336(.A (n_470), .B (n_196), .Y (n_171));
  NAND2X1 g1340(.A (n_150), .B (n_128), .Y (n_194));
  NAND2X1 g1343(.A (rtr), .B (n_460), .Y (n_377));
  AND2X1 g1345(.A (n_190), .B (n_381), .Y (n_207));
  NAND2X1 g1346(.A (n_148), .B (n_215), .Y (n_169));
  NAND3X1 g1348(.A (n_409), .B (start), .C (n_154), .Y (n_168));
  NAND3X1 g1350(.A (n_406), .B (n_178), .C (n_1), .Y (n_167));
  NAND2X1 g1351(.A (n_148), .B (n_190), .Y (n_166));
  NAND3X1 g1353(.A (n_406), .B (start), .C (n_163), .Y (n_165));
  NAND2X1 g1355(.A (n_85), .B (n_460), .Y (n_162));
  CLKBUFX3 g1385(.A (n_191), .Y (n_223));
  INVX2 g1399(.A (n_388), .Y (n_251));
  INVX1 g1402(.A (n_389), .Y (n_186));
  NAND2X1 g1287(.A (n_182), .B (n_148), .Y (n_156));
  OAI21X1 g1239(.A0 (rtr), .A1 (n_154), .B0 (n_188), .Y (n_155));
  INVX1 g1330(.A (n_182), .Y (n_153));
  NAND2X1 g1333(.A (n_135), .B (n_163), .Y (n_152));
  NAND2X1 g1337(.A (n_135), .B (n_150), .Y (n_151));
  INVX1 g1362(.A (n_230), .Y (n_149));
  INVX1 g1367(.A (n_175), .Y (n_161));
  INVX2 g1374(.A (n_148), .Y (n_249));
  INVX1 g1380(.A (n_460), .Y (n_145));
  INVX4 g1388(.A (n_142), .Y (n_191));
  INVX1 g1392(.A (n_381), .Y (n_204));
  INVX1 g1396(.A (n_406), .Y (n_141));
  CLKBUFX3 g1405(.A (n_431), .Y (n_221));
  NAND4X1 g1282(.A (rtr), .B (n_72), .C (n_137), .D (n_348), .Y
       (n_138));
  NAND3X1 g1331(.A (n_1), .B (n_137), .C (n_125), .Y (n_182));
  INVX2 g1368(.A (n_133), .Y (n_175));
  INVX2 g1358(.A (n_132), .Y (n_256));
  INVX1 g1359(.A (n_132), .Y (n_131));
  INVX2 g1363(.A (n_449), .Y (n_230));
  CLKBUFX3 g1364(.A (n_449), .Y (n_215));
  INVX2 g1376(.A (n_135), .Y (n_148));
  INVX2 g1389(.A (n_123), .Y (n_142));
  CLKBUFX3 g1407(.A (n_190), .Y (n_196));
  INVX1 g1408(.A (n_190), .Y (n_128));
  NAND2X1 g1283(.A (n_87), .B (key), .Y (n_127));
  NAND3X1 g1284(.A (n_104), .B (n_391), .C (n_125), .Y (n_126));
  NAND2X1 g1286(.A (n_98), .B (key), .Y (n_124));
  NAND2X2 g1390(.A (n_122), .B (n_113), .Y (n_123));
  MX2X1 g1307(.A (n_300), .B (n_60), .S0 (start), .Y (n_121));
  MX2X1 g1308(.A (n_38), .B (n_67), .S0 (start), .Y (n_120));
  NAND3X1 g1316(.A (rts), .B (n_122), .C (n_348), .Y (n_294));
  NAND2X1 g1252(.A (n_77), .B (rtr), .Y (n_188));
  NAND2X1 g1369(.A (n_137), .B (n_125), .Y (n_133));
  INVX2 g1377(.A (n_115), .Y (n_135));
  INVX1 g1360(.A (n_97), .Y (n_132));
  NAND2X2 g1409(.A (n_137), .B (n_113), .Y (n_190));
  XOR2X1 g1276(.A (n_47), .B (n_63), .Y (n_112));
  OR2X1 g1424(.A (rtr), .B (n_99), .Y (n_111));
  INVX2 g1425(.A (n_110), .Y (n_140));
  NAND2X1 g1378(.A (n_404), .B (n_456), .Y (n_115));
  NOR2X1 g1321(.A (n_103), .B (n_73), .Y (n_104));
  XOR2X1 g1357(.A (n_79), .B (n_34), .Y (n_98));
  NAND2X1 g1361(.A (n_122), .B (n_125), .Y (n_97));
  MX2X1 g1412(.A (n_4), .B (n_15), .S0 (rtr), .Y (n_96));
  MX2X1 g1413(.A (n_2), .B (n_31), .S0 (rtr), .Y (n_95));
  OAI21X1 g1414(.A0 (rts), .A1 (n_15), .B0 (n_16), .Y (n_94));
  MX2X1 g1415(.A (n_5), .B (n_61), .S0 (rtr), .Y (n_92));
  OAI21X1 g1416(.A0 (n_15), .A1 (start), .B0 (n_29), .Y (n_91));
  OAI21X1 g1418(.A0 (rts), .A1 (n_61), .B0 (n_13), .Y (n_90));
  OAI21X1 g1419(.A0 (n_246), .A1 (n_31), .B0 (n_8), .Y (n_89));
  INVX2 g1426(.A (n_402), .Y (n_110));
  XOR2X1 g1356(.A (n_61), .B (n_36), .Y (n_87));
  NAND2X1 g1455(.A (n_1), .B (n_49), .Y (n_86));
  NAND2X1 g1431(.A (rtr), .B (n_74), .Y (n_85));
  OAI21X1 g1411(.A0 (rts), .A1 (n_79), .B0 (n_22), .Y (n_80));
  MX2X1 g1420(.A (n_7), .B (n_79), .S0 (rtr), .Y (n_78));
  NAND3X1 g1280(.A (n_30), .B (n_15), .C (n_31), .Y (n_77));
  INVX2 g1432(.A (n_454), .Y (n_137));
  INVX2 g1435(.A (n_57), .Y (n_113));
  OR2X1 g1439(.A (rtr), .B (n_74), .Y (n_75));
  INVX1 g1473(.A (n_72), .Y (n_99));
  NOR2X1 g1410(.A (n_24), .B (n_21), .Y (n_103));
  INVX1 g1527(.A (n_61), .Y (n_244));
  OAI21X1 g1417(.A0 (n_33), .A1 (key), .B0 (n_17), .Y (n_67));
  INVX1 g1474(.A (n_73), .Y (n_72));
  INVX1 g1509(.A (n_74), .Y (n_163));
  XOR2X1 g1422(.A (n_79), .B (n_61), .Y (n_63));
  OAI21X1 g1421(.A0 (n_35), .A1 (key), .B0 (n_12), .Y (n_60));
  NOR2X1 g1423(.A (n_79), .B (start), .Y (n_59));
  INVX1 g1457(.A (n_403), .Y (n_122));
  NAND2X2 g1436(.A (n_39), .B (n_37), .Y (n_57));
  INVX2 g1450(.A (n_447), .Y (n_125));
  INVX1 g1496(.A (n_154), .Y (n_470));
  INVX1 g1513(.A (n_269), .Y (n_49));
  INVX1 g1475(.A (n_465), .Y (n_73));
  INVX1 g1498(.A (n_462), .Y (n_350));
  INVX1 g1514(.A (n_39), .Y (n_269));
  INVX1 g1510(.A (n_37), .Y (n_74));
  NAND2X1 g1438(.A (n_35), .B (g_button), .Y (n_36));
  NAND2X1 g1437(.A (n_33), .B (r_button), .Y (n_34));
  NOR2X1 g1453(.A (n_79), .B (n_61), .Y (n_30));
  NAND2X1 g1454(.A (key), .B (start), .Y (n_29));
  CLKBUFX1 g1497(.A (n_462), .Y (n_154));
  NAND2X1 g1460(.A (v_in[0]), .B (v_in[1]), .Y (n_24));
  INVX1 g1518(.A (n_150), .Y (n_246));
  NAND2X1 g1443(.A (v_in[2]), .B (rts), .Y (n_22));
  NAND2X1 g1445(.A (v_in[2]), .B (v_in[3]), .Y (n_21));
  NOR2X1 g1461(.A (rtr), .B (cts), .Y (n_20));
  INVX1 g1511(.A (n_46), .Y (n_37));
  NAND2X1 g1456(.A (r_button), .B (key), .Y (n_17));
  NAND2X1 g1449(.A (v_in[0]), .B (rts), .Y (n_16));
  NAND2X1 g1442(.A (v_in[1]), .B (rts), .Y (n_13));
  NAND2X1 g1447(.A (g_button), .B (key), .Y (n_12));
  INVX2 g1516(.A (n_45), .Y (n_9));
  NAND2X1 g1446(.A (rts), .B (v_in[3]), .Y (n_8));
  CLKBUFX2 g1515(.A (n_45), .Y (n_39));
  INVX1 g1526(.A (n_47), .Y (n_15));
  INVX1 g1485(.A (v_out[2]), .Y (n_7));
  INVX1 g1502(.A (n_300), .Y (n_35));
  INVX4 g1512(.A (stato_6), .Y (n_46));
  INVX1 g1520(.A (rts), .Y (n_150));
  INVX1 g1482(.A (v_in[3]), .Y (n_6));
  INVX1 g1521(.A (reset), .Y (n_340));
  INVX1 g1484(.A (v_out[1]), .Y (n_5));
  INVX1 g1478(.A (v_out[0]), .Y (n_4));
  INVX1 g1467(.A (n_27), .Y (n_31));
  INVX2 g1517(.A (stato_5), .Y (n_45));
  INVX1 g1483(.A (v_out[3]), .Y (n_2));
  INVX1 g1531(.A (n_178), .Y (n_61));
  INVX1 g1491(.A (start), .Y (n_1));
  INVX1 g1506(.A (n_286), .Y (n_18));
  INVX1 g1481(.A (n_38), .Y (n_33));
  INVX2 g1535(.A (voto2), .Y (n_79));
  CLKBUFX1 g1554(.A (n_456), .Y (n_348));
  NAND2X1 g1393_dup(.A (n_451), .B (n_125), .Y (n_381));
  NAND2X2 g1574(.A (n_140), .B (n_137), .Y (n_388));
  NAND2X2 g1403_dup(.A (n_140), .B (n_137), .Y (n_389));
  NOR2X1 g1575(.A (n_350), .B (n_73), .Y (n_466));
  NOR2X1 g1448_dup(.A (n_350), .B (n_73), .Y (n_391));
  INVX1 g1576(.A (n_453), .Y (n_392));
  AND2X1 g41(.A (n_400), .B (n_407), .Y (n_408));
  NAND2X1 g42(.A (n_397), .B (n_399), .Y (n_400));
  NAND3X1 g43(.A (n_27), .B (start), .C (key), .Y (n_397));
  INVX1 g47(.A (n_398), .Y (n_399));
  NOR2X1 g48(.A (start), .B (n_31), .Y (n_398));
  CLKBUFX3 g53(.A (n_406), .Y (n_407));
  INVX2 g54(.A (n_405), .Y (n_406));
  NAND2X1 g46(.A (n_402), .B (n_404), .Y (n_405));
  INVX2 g51(.A (n_401), .Y (n_402));
  NAND2X2 g52(.A (n_9), .B (n_46), .Y (n_401));
  INVX1 g49(.A (n_403), .Y (n_404));
  NAND2X1 g50(.A (n_461), .B (n_463), .Y (n_403));
  CLKBUFX2 g1(.A (n_406), .Y (n_409));
  NAND4X1 g1579(.A (n_411), .B (n_412), .C (n_413), .D (n_415), .Y
       (n_416));
  AOI21X1 g44(.A0 (ctr), .A1 (n_459), .B0 (n_195), .Y (n_411));
  OAI21X1 g45(.A0 (n_287), .A1 (n_407), .B0 (ctr), .Y (n_412));
  NAND2X1 g1581(.A (n_197), .B (ctr), .Y (n_413));
  NAND2X1 g1582(.A (n_414), .B (ctr), .Y (n_415));
  NAND3X1 g1583(.A (n_151), .B (n_215), .C (n_432), .Y (n_414));
  NAND2X1 g17(.A (n_430), .B (n_432), .Y (n_433));
  NAND2X1 g18(.A (rtr), .B (n_459), .Y (n_430));
  INVX2 g19(.A (n_431), .Y (n_432));
  NOR2X1 g20(.A (n_464), .B (n_110), .Y (n_431));
  NAND2X2 g36(.A (n_444), .B (n_445), .Y (n_446));
  NOR2X1 g37(.A (n_442), .B (n_443), .Y (n_444));
  OAI21X1 g38(.A0 (n_441), .A1 (n_381), .B0 (n_200), .Y (n_442));
  AND2X1 g1596(.A (n_99), .B (rtr), .Y (n_441));
  NAND3X1 g39(.A (n_241), .B (n_218), .C (n_294), .Y (n_443));
  AOI21X1 g40(.A0 (n_174), .A1 (n_246), .B0 (n_214), .Y (n_445));
  NAND2X1 g1597(.A (n_449), .B (n_458), .Y (n_453));
  NAND2X2 g1598(.A (n_125), .B (n_466), .Y (n_449));
  NAND2X1 g26(.A (n_46), .B (n_45), .Y (n_447));
  INVX1 g1599(.A (n_464), .Y (n_451));
  NAND2X1 g1601(.A (n_457), .B (n_458), .Y (n_459));
  NAND2X2 g1602(.A (n_455), .B (n_456), .Y (n_457));
  INVX1 g28(.A (n_454), .Y (n_455));
  NAND2X2 g29(.A (n_465), .B (n_461), .Y (n_454));
  NOR2X1 g30(.A (n_45), .B (n_46), .Y (n_456));
  NAND2X1 g27(.A (n_451), .B (n_125), .Y (n_458));
  INVX2 g1603(.A (n_457), .Y (n_460));
  NAND2X1 g11(.A (n_462), .B (n_463), .Y (n_464));
  INVX1 g14(.A (n_461), .Y (n_462));
  INVX2 g15(.A (stato_7), .Y (n_461));
  INVX2 g13(.A (stato), .Y (n_463));
  INVX2 g12(.A (n_463), .Y (n_465));
endmodule

