//
//  ITC99 Benchmark
//  Downloaded from http://www.cad.polito.it/tools/itc99.html
//  
//  ----------------------------------------------------------------------
//  
//  This netlist was generated with Cadence RTL Compiler in a quick 
//  synthesis run.
//  
//  ----------------------------------------------------------------------
//  
//  Copyright (C) 1999
//  Fulvio Corno, Matteo Sonze Reorda, Giovanni Squillero
//  Politecnico di Torino
//  
//  This source file may be used and distributed without restriction
//  provided that this copyright statement is not removed from the
//  file and that any derivative work contains the original copyright
//  notice and the associated disclaimer.
//  
//  This source file is free software; you can redistribute it and/or
//  modify it under the terms of the GNU General Public License as
//  published by the Free Software Foundation.
//  
//  This source is distributed in the hope that it will be useful,
//  but WITHOUT ANY WARRANTY; without even the implied warranty of
//  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
//  General Public License for more details.
//  
//  You should have received a copy of the GNU General Public License
//  along with this source; if not, download it from
//  http://www.gnu.org/copyleft/gpl.html
//  

// Generated by Cadence RTL Compiler (RC) v05.10-b006_1

module b06(cc_mux, eql, uscite, clock, enable_count, ackout, reset,
     cont_eql);
  input eql, clock, reset, cont_eql;
  output [2:1] cc_mux, uscite;
  output enable_count, ackout;
  wire eql, clock, reset, cont_eql;
  wire [2:1] cc_mux, uscite;
  wire enable_count, ackout;
  wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7;
  wire n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16;
  wire n_17, n_19, n_20, n_22, n_23, n_24, n_25, n_26;
  wire n_27, n_28, n_30, n_31, n_32, n_33, n_34, n_36;
  wire n_37, n_38, n_39, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53;
  wire n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69;
  wire n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77;
  wire n_78, n_79, n_80, n_83, n_84, state, state_7, state_8;
  DFFSRX1 \cc_mux_reg[1] (.RN (n_80), .SN (1'b1), .CK (clock), .D
       (n_78), .Q (cc_mux[1]), .QN ());
  DFFSRX1 enable_count_reg(.RN (n_80), .SN (1'b1), .CK (clock), .D
       (n_79), .Q (enable_count), .QN ());
  DFFSRX1 ackout_reg(.RN (n_80), .SN (1'b1), .CK (clock), .D (n_79), .Q
       (ackout), .QN ());
  DFFSRX1 \cc_mux_reg[2] (.RN (n_80), .SN (1'b1), .CK (clock), .D
       (n_77), .Q (cc_mux[2]), .QN ());
  DFFSRX1 \state_reg[1] (.RN (n_80), .SN (1'b1), .CK (clock), .D
       (n_76), .Q (state_7), .QN ());
  NAND2X2 g212(.A (n_74), .B (n_61), .Y (n_78));
  DFFSRX1 \state_reg[0] (.RN (n_80), .SN (1'b1), .CK (clock), .D
       (n_75), .Q (state), .QN ());
  DFFSRX1 \state_reg[2] (.RN (n_80), .SN (1'b1), .CK (clock), .D
       (n_73), .Q (state_8), .QN ());
  DFFSRX1 \uscite_reg[1] (.RN (n_80), .SN (1'b1), .CK (clock), .D
       (n_72), .Q (uscite[1]), .QN ());
  NAND2X2 g213(.A (n_69), .B (n_66), .Y (n_79));
  NAND2X2 g218(.A (n_67), .B (n_58), .Y (n_77));
  NAND2X2 g220(.A (n_71), .B (n_57), .Y (n_76));
  NAND3X1 g219(.A (n_62), .B (n_49), .C (n_31), .Y (n_75));
  INVX2 g215(.A (n_68), .Y (n_74));
  NAND3X1 g223(.A (n_64), .B (n_43), .C (n_31), .Y (n_73));
  NAND4X1 g211(.A (n_51), .B (n_37), .C (n_54), .D (n_46), .Y (n_72));
  NOR2X1 g225(.A (n_42), .B (n_70), .Y (n_71));
  DFFSRX1 \uscite_reg[2] (.RN (n_80), .SN (1'b1), .CK (clock), .D
       (n_70), .Q (uscite[2]), .QN ());
  NAND2X1 g222(.A (n_56), .B (n_65), .Y (n_69));
  NAND4X1 g216(.A (n_39), .B (n_41), .C (n_52), .D (n_45), .Y (n_68));
  NOR2X1 g224(.A (n_63), .B (n_44), .Y (n_67));
  AOI21X1 g217(.A0 (n_38), .A1 (n_65), .B0 (n_50), .Y (n_66));
  INVX1 g231(.A (n_63), .Y (n_64));
  NOR2X1 g234(.A (n_60), .B (n_53), .Y (n_62));
  NAND2X2 g227(.A (n_84), .B (n_59), .Y (n_70));
  NOR2X1 g230(.A (n_13), .B (n_60), .Y (n_61));
  NAND2X1 g232(.A (n_55), .B (n_59), .Y (n_63));
  AND2X1 g236(.A (n_47), .B (n_24), .Y (n_58));
  AOI21X1 g237(.A0 (n_36), .A1 (eql), .B0 (n_26), .Y (n_57));
  NAND4X1 g238(.A (n_55), .B (n_20), .C (n_33), .D (n_25), .Y (n_56));
  NOR2X1 g228(.A (n_48), .B (n_34), .Y (n_54));
  INVX1 g254(.A (n_52), .Y (n_53));
  NOR2X1 g229(.A (n_23), .B (n_50), .Y (n_51));
  NOR2X1 g235(.A (n_48), .B (n_50), .Y (n_49));
  NAND2X1 g244(.A (n_26), .B (eql), .Y (n_47));
  NOR2X1 g226(.A (n_19), .B (n_30), .Y (n_46));
  NAND2X1 g248(.A (n_27), .B (eql), .Y (n_45));
  INVX1 g249(.A (n_43), .Y (n_44));
  INVX1 g252(.A (n_41), .Y (n_42));
  NAND2X2 g255(.A (n_19), .B (n_1), .Y (n_52));
  NAND3X1 g233(.A (n_28), .B (n_24), .C (n_32), .Y (n_38));
  INVX1 g265(.A (n_36), .Y (n_37));
  NAND4X1 g239(.A (n_83), .B (n_16), .C (n_3), .D (eql), .Y (n_59));
  INVX1 g240(.A (n_34), .Y (n_84));
  NAND2X1 g242(.A (n_33), .B (n_32), .Y (n_60));
  INVX1 g245(.A (n_30), .Y (n_31));
  NAND2X1 g250(.A (n_14), .B (eql), .Y (n_43));
  NOR2X1 g251(.A (n_28), .B (eql), .Y (n_50));
  NAND2X1 g253(.A (n_17), .B (eql), .Y (n_41));
  INVX2 g258(.A (n_27), .Y (n_55));
  INVX1 g262(.A (n_26), .Y (n_39));
  INVX1 g266(.A (n_33), .Y (n_36));
  NOR2X1 g241(.A (n_22), .B (eql), .Y (n_34));
  NOR2X1 g243(.A (n_25), .B (eql), .Y (n_48));
  NOR2X1 g247(.A (n_24), .B (eql), .Y (n_30));
  INVX1 g256(.A (n_32), .Y (n_23));
  INVX2 g259(.A (n_22), .Y (n_27));
  INVX1 g263(.A (n_28), .Y (n_26));
  INVX2 g272(.A (n_20), .Y (n_19));
  NAND3X1 g267(.A (n_7), .B (n_16), .C (n_15), .Y (n_33));
  NAND3X1 g264(.A (n_16), .B (n_9), .C (n_15), .Y (n_28));
  NAND3X1 g260(.A (n_12), .B (n_10), .C (n_11), .Y (n_22));
  INVX1 g269(.A (n_25), .Y (n_14));
  INVX1 g268(.A (n_25), .Y (n_13));
  NAND3X1 g273(.A (n_12), .B (n_16), .C (n_11), .Y (n_20));
  NAND3X1 g257(.A (n_9), .B (n_10), .C (n_15), .Y (n_32));
  INVX1 g275(.A (n_24), .Y (n_17));
  NAND2X2 g270(.A (n_5), .B (n_10), .Y (n_25));
  NAND3X1 g276(.A (n_0), .B (n_6), .C (n_15), .Y (n_24));
  INVX1 g286(.A (n_7), .Y (n_83));
  INVX2 g287(.A (n_9), .Y (n_7));
  INVX2 g285(.A (n_6), .Y (n_12));
  NOR2X1 g277(.A (n_2), .B (n_4), .Y (n_5));
  INVX2 g288(.A (n_6), .Y (n_9));
  INVX1 g283(.A (n_4), .Y (n_11));
  INVX1 g281(.A (n_15), .Y (n_3));
  INVX4 g289(.A (n_2), .Y (n_6));
  INVX1 g278(.A (reset), .Y (n_80));
  INVX1 g279(.A (eql), .Y (n_1));
  INVX1 g292(.A (state_7), .Y (n_0));
  INVX1 g284(.A (state_8), .Y (n_4));
  INVX1 g291(.A (state_7), .Y (n_10));
  INVX1 g282(.A (state_8), .Y (n_15));
  INVX2 g290(.A (state), .Y (n_2));
  INVX1 g280(.A (cont_eql), .Y (n_65));
  CLKBUFX1 g293(.A (state_7), .Y (n_16));
endmodule

